--controls the entire operation
--via control signals taken from stage units and driven to later stage ones
--and enable signals of input and output regs

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity control_unit is
	port(--clock and reset input signals
	     clk,rst: in std_logic;

	     --signal to start the operations
	     start: in std_logic;
	     
	     --control input signals
	     spec_case: in std_logic;                          --initial input special case check
	     cmp: in std_logic;                                --exponent compare
	     shift_num: in std_logic_vector(4 downto 0);       --number of shifts needed in mantissa
	     cout: in std_logic;                               --carry out from mantissa addition
	     round_ovf: in std_logic;                          --overflow in rounding
	     inc_dec_inf: in std_logic;                        --infinity in increament/decreament of exponent
             inc_dec_unf: in std_logic;                        --underflow in increament/decreament of exponent
	     
	     --output control signals
	     out_flags: out std_logic_vector(10 downto 0);     --control flags needed in different units
	     regs_control: out std_logic_vector(3 downto 0)    --inreg_wr & inreg_rd & outreg_wr & outreg_rd

	     --done: out std_logic;
	    );
end control_unit;
architecture control_unit_arch of control_unit is 

--states declaration
type state is (wait_state, yellow_state, rose_state, red_state, lblue_state, dblue_state);
signal pr_state, nx_state: state;

--mid signals
signal mid_flags: std_logic_vector(10 downto 0);
begin
	mid_flags <= spec_case & cmp & shift_num & cout & round_ovf & inc_dec_inf & inc_dec_unf;
	out_flags <= mid_flags;
	
	--clock and reset process
	P1: process(clk,rst)
	begin
		if(rst='1') then
			pr_state <= wait_state;
		elsif(clk'event and clk='1') then
			pr_state <= nx_state;
		end if;
	end process P1;

	--next state and output process
	P2: process(spec_case,pr_state)   -----or mid_flags?
	begin
		case pr_state is
			when wait_state => 
				regs_control <= "1000";
				out_flags <= "XXXXXXXXXXX";
				if(start='1') then  
					nx_state <= yellow_state;
				else
					nx_state <= wait_state;
				end if;
			when yellow_state =>
				regs_control <= "0100";
				if(spec_case='1') then   -----or mid_flags?
					nx_state <= rose_state;
				else
					nx_state <= dblue_state;
				end if;
			when rose_state =>
				regs_control <= "0000";
				nx_state <= red_state;
			when red_state =>
				regs_control <= "0000";
				nx_state <= lblue_state;
			when lblue_state => 
				regs_control <= "0000";
				nx_state <= dblue_state;
			when dblue_state =>
				regs_control <= "0011"; ----????
				nx_state <= wait_state;
		end case;
	end process P2;
end control_unit_arch;
