--register that stores the sum output of the fp adder and its flags

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity output_register is
	port(clk,rst: in std_logic;
	     wr_en: in std_logic;
	     sum_in: in std_logic_vector(31 downto 0);        --the sum of the fp adder
             unf_flag_in: in std_logic;                       --underflow flag in the case where the exponent after the inc/dec stage becomes zero
	     sum_out: out std_logic_vector(31 downto 0);
             unf_flag_out: out std_logic
	     );
end output_register;

architecture output_register_arch of output_register is
	signal reg: std_logic_vector(31 downto 0);
	signal unf_flag: std_logic;
begin
	process(clk,rst)
        begin
        	if(rst = '1') then
                	reg <= (others =>'0');
			unf_flag <= '0';
                elsif(clk'event and clk = '1') then                         
                	if(wr_en = '1') then
                		reg <= sum_in;
				unf_flag <= unf_flag_in;
                        end if;
                end if;
        end process;
	
	sum_out <= reg;                                              
	unf_flag_out <= unf_flag;
		       
end output_register_arch;
